//-----
// Parse Data Signal for bits
//-----
// ensure ps2_data bit[0] = 0

// parse ps2_data bit[1:8] for actual data

// examine ps2_data bit[9] as odd parity bit; ensure data is correct.

// ensure ps2_data bit[10] = 1

